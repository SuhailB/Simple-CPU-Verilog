//module MAR(clk, reset, write, read, in_from_bus, out_to_bus); //read is not necessary
module MAR  (clk, reset, in_from_bus, out_to_bus, write, mem_read); 

input clk, reset, write, read;
input [15:0] in_from_bus;
output[15:0] out_to_bus;

reg[15:0] register;

always@(posedge clk or posedge reset)
begin
  if(reset) register <= 0;
  else if(write) register <= in_from_bus;
end

assign out_to_bus = mem_read? register : 16'hzzzz;

endmodule